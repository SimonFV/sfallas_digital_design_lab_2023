module check_defeat();


endmodule