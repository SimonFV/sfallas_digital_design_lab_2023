module main(output logic pc);

	assign pc = 1;

endmodule