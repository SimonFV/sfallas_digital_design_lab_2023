module color(input int value, output [23:0] pixel_color);
	
	always_comb begin
		case (value)
			0: pixel_color = 24'b000111000001110000011100;
			2: pixel_color = 24'b111111111111111111001100;
			4: pixel_color = 24'b111111111111111111100110;
			8: pixel_color = 24'b111111111100110010011001;
			16: pixel_color = 24'b111111111100110011001100;
			32: pixel_color = 24'b111111111100110010011001;
			64: pixel_color = 24'b111111111001100110011001;
			128: pixel_color = 24'b111111111100110011001100;
			256: pixel_color = 24'b111111111001100111001100;
			512: pixel_color = 24'b110011000110011001100110;
			1024: pixel_color = 24'b100110010011001100110011;
			2048: pixel_color = 24'b110011001111111111001100;
			100: pixel_color = 24'b000011000000110000001100;
			default: pixel_color = 24'b000011000000110000001100;
		endcase
	end
	
endmodule