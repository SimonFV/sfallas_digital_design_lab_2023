module color(input [3:0] value, output [23:0] pixel_color);
	
	always_comb begin
		case (value)
			0: pixel_color = 24'b111111111111111110011001;
			1: pixel_color = 24'b111111111111111111001100;
			2: pixel_color = 24'b111111111111111111100110;
			3: pixel_color = 24'b111111111100110010011001;
			4: pixel_color = 24'b111111111100110011001100;
			5: pixel_color = 24'b111111111100110010011001;
			6: pixel_color = 24'b111111111001100110011001;
			7: pixel_color = 24'b111111111100110011001100;
			8: pixel_color = 24'b111111111001100111001100;
			9: pixel_color = 24'b110011000110011001100110;
			10: pixel_color = 24'b100110010011001100110011;
			11: pixel_color = 24'b110011001111111111001100;
			default: pixel_color = 24'b110111001101110011011100;
		endcase
	end
	
endmodule