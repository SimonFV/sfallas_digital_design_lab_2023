module alu_not (input logic a, output logic result);

assign result = ~a;

endmodule
