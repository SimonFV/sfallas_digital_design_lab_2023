module decodificador();


endmodule
