module color(input [3:0] value, output [23:0] pixel_color);
	
	always_comb begin
		case (value)
			4'b0000: pixel_color = 24'b111111111111111110011001;
			4'b0001: pixel_color = 24'b111111111111111111001100;
			4'b0010: pixel_color = 24'b111111111111111111100110;
			4'b0011: pixel_color = 24'b111111111100110010011001;
			4'b0100: pixel_color = 24'b111111111100110011001100;
			4'b0101: pixel_color = 24'b111111111100110010011001;
			4'b0110: pixel_color = 24'b111111111001100110011001;
			4'b0111: pixel_color = 24'b111111111100110011001100;
			4'b1000: pixel_color = 24'b111111111001100111001100;
			4'b1001: pixel_color = 24'b110011000110011001100110;
			4'b1010: pixel_color = 24'b100110010011001100110011;
			4'b1011: pixel_color = 24'b110011001111111111001100;
			default: pixel_color = 24'b110111001101110011011100;
		endcase
	end
	
endmodule